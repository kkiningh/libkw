`default_nettype none

module SRAM1RW32x50 (
  input wire [5-1:0] A,
  input wire CE,
  input wire WEB,
  input wire OEB,
  input wire CSB,
  input wire [50-1:0] I,
  output reg [50-1:0] O
);
  wire RE = ~CSB && WEB;
  wire WE = ~CSB && ~WEB;

  reg [32-1:0][50-1:0] mem;
  reg [50-1:0] data_out;
  always_ff @(posedge CE) begin
    if (RE) data_out <= mem[A];
    if (WE) mem[A] <= I;
  end

  assign O = !OEB ? data_out : 50'bz;
endmodule
