`default_nettype none

/* verilator lint_off UNUSED */
module KW_unread (
  input logic d_i
);

endmodule
/* verilator lint_on UNUSED */
